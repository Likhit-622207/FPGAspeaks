module not_1(
    input a,
    output b
    );
assign b=~a;
endmodule
