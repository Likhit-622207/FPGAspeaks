 module and_2(
    input a,b,
    output c
    );
    assign c=a&b;
endmodule
